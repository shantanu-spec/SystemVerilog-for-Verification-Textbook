//Given Binary::copy function create ExtBinary copy
class Binary;
  rand bit [3:0] val1, val2;
  
  function new(input bit [3:0] val1,val2);
		this.val1 = val1;
    	this.val2 = val2;
  endfunction: new
  
  virtual function void print_int(input int val);
    $display("val=0d%0d",val);
  endfunction: print_int
  
  virtual function Binary copy();
    copy = new(15,8);
    copy.val1 = val1;
  	copy.val2 = val2;
  endfunction: copy
  
endclass: Binary

class ExtBinary extends Binary;
  
  function new(input bit [3:0] val1,val2);
    super.new(val1,val2);
  endfunction: new
  
  virtual function int mult_val();
    return val1*val2;
  endfunction:mult_val
  
  virtual function Binary copy();
  	ExtBinary copy;
  	copy = new(this.val1, this.val2); 
    return copy;
  endfunction: copy
  
endclass: ExtBinary

class Exercise3 extends ExtBinary;
  
  function new(input bit [3:0] val1,val2);
    super.new(val1,val2);
  endfunction: new
  
  constraint val1set {val1 < 10;}
  constraint val2set {val2 < 10;}
endclass: Exercise3

module ex3;
  Exercise3 ex3;
  initial begin
    
    ex3 = new(0,0);
    if(!ex3.randomize())
      $display("Randomization ERROR!");
    else
      ex3.print_int(ex3.val1);
      ex3.print_int(ex3.val2);
      ex3.print_int(ex3.mult_val());
    
  end
endmodule
